module verificador_paridade_tb;
    
    reg b1, b2, b3, b4, b5, bp; //entradas
    wire S; //saida          

    verificador_paridade teste(  
        .b1(b1), //faz a conexão com o modulo
        .b2(b2),
        .b3(b3),
        .b4(b4),
        .b5(b5),
        .bp(bp),
        .S(S)
    );

    initial begin

        $display("b1 b2 b3 b4 b5 bp - S");
        $monitor("%b  %b  %b  %b  %b  %b  %b", b1, b2, b3, b4, b5, bp, S);

        b1= 0; b2= 0; b3= 0; b4= 0; b5= 0; bp= 0;#10; //tabela verdade
        b1= 0; b2= 0; b3= 0; b4= 0; b5= 0; bp= 1;#10; //obs, verificar se esse tempo de atraso é suficiente
        b1= 0; b2= 0; b3= 0; b4= 0; b5= 1; bp= 0;#10; 
        b1= 0; b2= 0; b3= 0; b4= 0; b5= 1; bp= 1;#10; 
        b1= 0; b2= 0; b3= 0; b4= 1; b5= 0; bp= 0;#10; 
        b1= 0; b2= 0; b3= 0; b4= 1; b5= 0; bp= 1;#10; 
        b1= 0; b2= 0; b3= 0; b4= 1; b5= 1; bp= 0;#10; 
        b1= 0; b2= 0; b3= 0; b4= 1; b5= 1; bp= 1;#10; 
        b1= 0; b2= 0; b3= 1; b4= 0; b5= 0; bp= 0;#10; 
        b1= 0; b2= 0; b3= 1; b4= 0; b5= 0; bp= 1;#10; 
        b1= 0; b2= 0; b3= 1; b4= 0; b5= 1; bp= 0;#10; 
        b1= 0; b2= 0; b3= 1; b4= 0; b5= 1; bp= 1;#10; 
        b1= 0; b2= 0; b3= 1; b4= 1; b5= 0; bp= 0;#10; 
        b1= 0; b2= 0; b3= 1; b4= 1; b5= 0; bp= 1;#10; 
        b1= 0; b2= 0; b3= 1; b4= 1; b5= 1; bp= 0;#10; 
        b1= 0; b2= 0; b3= 1; b4= 1; b5= 1; bp= 1;#10; 

        b1= 0; b2= 1; b3= 0; b4= 0; b5= 0; bp= 0;#10;
        b1= 0; b2= 1; b3= 0; b4= 0; b5= 0; bp= 1;#10;
        b1= 0; b2= 1; b3= 0; b4= 0; b5= 1; bp= 0;#10;
        b1= 0; b2= 1; b3= 0; b4= 0; b5= 1; bp= 1;#10; 
        b1= 0; b2= 1; b3= 0; b4= 1; b5= 0; bp= 0;#10; 
        b1= 0; b2= 1; b3= 0; b4= 1; b5= 0; bp= 1;#10;
        b1= 0; b2= 1; b3= 0; b4= 1; b5= 1; bp= 0;#10;
        b1= 0; b2= 1; b3= 0; b4= 1; b5= 1; bp= 1;#10;
        b1= 0; b2= 1; b3= 1; b4= 0; b5= 0; bp= 0;#10;
        b1= 0; b2= 1; b3= 1; b4= 0; b5= 0; bp= 1;#10;
        b1= 0; b2= 1; b3= 1; b4= 0; b5= 1; bp= 0;#10;
        b1= 0; b2= 1; b3= 1; b4= 0; b5= 1; bp= 1;#10;
        b1= 0; b2= 1; b3= 1; b4= 1; b5= 0; bp= 0;#10;
        b1= 0; b2= 1; b3= 1; b4= 1; b5= 0; bp= 1;#10;
        b1= 0; b2= 1; b3= 1; b4= 1; b5= 1; bp= 0;#10;
        b1= 0; b2= 1; b3= 1; b4= 1; b5= 1; bp= 1;#10;

        b1= 1; b2= 0; b3= 0; b4= 0; b5= 0; bp= 0;#10;
        b1= 1; b2= 0; b3= 0; b4= 0; b5= 0; bp= 1;#10;
        b1= 1; b2= 0; b3= 0; b4= 0; b5= 1; bp= 0;#10;
        b1= 1; b2= 0; b3= 0; b4= 0; b5= 1; bp= 1;#10;
        b1= 1; b2= 0; b3= 0; b4= 1; b5= 0; bp= 0;#10;
        b1= 1; b2= 0; b3= 0; b4= 1; b5= 0; bp= 1;#10;
        b1= 1; b2= 0; b3= 0; b4= 1; b5= 1; bp= 0;#10;
        b1= 1; b2= 0; b3= 0; b4= 1; b5= 1; bp= 1;#10;
        b1= 1; b2= 0; b3= 1; b4= 0; b5= 0; bp= 0;#10;
        b1= 1; b2= 0; b3= 1; b4= 0; b5= 0; bp= 1;#10;
        b1= 1; b2= 0; b3= 1; b4= 0; b5= 1; bp= 0;#10;
        b1= 1; b2= 0; b3= 1; b4= 0; b5= 1; bp= 1;#10;
        b1= 1; b2= 0; b3= 1; b4= 1; b5= 0; bp= 0;#10;
        b1= 1; b2= 0; b3= 1; b4= 1; b5= 0; bp= 1;#10;
        b1= 1; b2= 0; b3= 1; b4= 1; b5= 1; bp= 0;#10;
        b1= 1; b2= 0; b3= 1; b4= 1; b5= 1; bp= 1;#10;

        b1= 1; b2= 1; b3= 0; b4= 0; b5= 0; bp= 0;#10;
        b1= 1; b2= 1; b3= 0; b4= 0; b5= 0; bp= 1;#10;
        b1= 1; b2= 1; b3= 0; b4= 0; b5= 1; bp= 0;#10;
        b1= 1; b2= 1; b3= 0; b4= 0; b5= 1; bp= 1;#10;
        b1= 1; b2= 1; b3= 0; b4= 1; b5= 0; bp= 0;#10;
        b1= 1; b2= 1; b3= 0; b4= 1; b5= 0; bp= 1;#10;
        b1= 1; b2= 1; b3= 0; b4= 1; b5= 1; bp= 0;#10;
        b1= 1; b2= 1; b3= 0; b4= 1; b5= 1; bp= 1;#10;
        b1= 1; b2= 1; b3= 1; b4= 0; b5= 0; bp= 0;#10;
        b1= 1; b2= 1; b3= 1; b4= 0; b5= 0; bp= 1;#10;
        b1= 1; b2= 1; b3= 1; b4= 0; b5= 1; bp= 0;#10;
        b1= 1; b2= 1; b3= 1; b4= 0; b5= 1; bp= 1;#10;
        b1= 1; b2= 1; b3= 1; b4= 1; b5= 0; bp= 0;#10;
        b1= 1; b2= 1; b3= 1; b4= 1; b5= 0; bp= 1;#10;
        b1= 1; b2= 1; b3= 1; b4= 1; b5= 1; bp= 0;#10;
        b1= 1; b2= 1; b3= 1; b4= 1; b5= 1; bp= 1;#10;


        $finish; 
    end
endmodule
