module display-7_seg (b1,b2,b3,b4,b5,b_par,A,B,C,D,E,F,G);
    input b1,b2,b3,b4,b5,b_par;
    output reg A,B,C,D,E,F,G;

    always@(*) begin
        if
        A <=
    end
endmodule